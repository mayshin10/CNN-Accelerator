`timescale 1ps / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/11/11 17:24:07
// Design Name: 
// Module Name: test_bench
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module test_bench();
    reg clk;
    reg reset;
    wire [31:0] AHB_INTERFACE_0_haddr;
    wire [2:0] AHB_INTERFACE_0_hburst;
    wire [3:0] AHB_INTERFACE_0_hprot;
    reg [31:0] AHB_INTERFACE_0_hrdata;
    wire AHB_INTERFACE_0_hready_in;
    reg AHB_INTERFACE_0_hready_out;
    reg AHB_INTERFACE_0_hresp;
    wire [2:0] AHB_INTERFACE_0_hsize;
    wire [1:0] AHB_INTERFACE_0_htrans;
    wire [31:0] AHB_INTERFACE_0_hwdata;
    wire AHB_INTERFACE_0_hwrite;
    wire AHB_INTERFACE_0_sel;
    reg start;
    wire finish;
    wire state_test;

    
   
    
    vector_add sim(
    .clk(clk),
    .reset(reset),
    .AHB_INTERFACE_0_haddr(AHB_INTERFACE_0_haddr),
        .AHB_INTERFACE_0_hburst(AHB_INTERFACE_0_hburst),
        .AHB_INTERFACE_0_hprot(AHB_INTERFACE_0_hprot),
        .AHB_INTERFACE_0_hrdata(AHB_INTERFACE_0_hrdata),
        .AHB_INTERFACE_0_hready_in(AHB_INTERFACE_0_hready_in),
        .AHB_INTERFACE_0_hready_out(AHB_INTERFACE_0_hready_out),
        .AHB_INTERFACE_0_hresp(AHB_INTERFACE_0_hresp),
        .AHB_INTERFACE_0_hsize(AHB_INTERFACE_0_hsize),
        .AHB_INTERFACE_0_htrans(AHB_INTERFACE_0_htrans),
        .AHB_INTERFACE_0_hwdata(AHB_INTERFACE_0_hwdata),
        .AHB_INTERFACE_0_hwrite(AHB_INTERFACE_0_hwrite),
        .AHB_INTERFACE_0_sel(AHB_INTERFACE_0_sel),
        .start(start),
        .finish(finish),
        .state_test(state_test)
        );

        initial begin
            clk <= 1'b0;
            reset <= 1'b0;
            AHB_INTERFACE_0_hready_out <=1'b1;
            AHB_INTERFACE_0_hresp<= 1'b0;
            #30
            reset <= 1'b1;
            start<=1;
         end
         always@(*)
         begin
         #10 clk <= ~clk;
            case(AHB_INTERFACE_0_haddr)//address_offset 확인 
         (32'h4001_0000+0): begin 
          AHB_INTERFACE_0_hrdata<=32'hd132ec2e; 
          end
         (32'h4001_0000+4): begin 
          AHB_INTERFACE_0_hrdata<=32'hf5efeb1f; 
          end
         (32'h4001_0000+8): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000025; 
          end
          (32'h4000_0000+0): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+8): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+12): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+16): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+20): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+24): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+28): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+32): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+36): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+40): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+44): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+48): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+52): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+56): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+60): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+64): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+68): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+72): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+76): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+80): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+84): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+88): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+92): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+96): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+100): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+104): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+108): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+112): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+116): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+120): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+124): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+128): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+132): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+136): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+140): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+144): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+148): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+152): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+156): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+160): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+164): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+168): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+172): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+176): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+180): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+184): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+188): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+192): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+196): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+200): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+204): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+208): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+212): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+216): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+220): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+224): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+228): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+232): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+236): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+240): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+244): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+248): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+252): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+256): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+260): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+264): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+268): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+272): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+276): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+280): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+284): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+288): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+292): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+296): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+300): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+304): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+308): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+312): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+316): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+320): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+324): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+328): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+332): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+336): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+340): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+344): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+348): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+352): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+356): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+360): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+364): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+368): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+372): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+376): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+380): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+384): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+388): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+392): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+396): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+400): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+404): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+408): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+412): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+416): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+420): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+424): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+428): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+432): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+436): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+440): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+444): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+448): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+452): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+456): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+460): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+464): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+468): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+472): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+476): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+480): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+484): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+488): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+492): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+496): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+500): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+504): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+508): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+512): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+516): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+520): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+524): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+528): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+532): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+536): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+540): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+544): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+548): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+552): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+556): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+560): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+564): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+568): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+572): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+576): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+580): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+584): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+588): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+592): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+596): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+600): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+604): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+608): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+612): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+616): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+620): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+624): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+628): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+632): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+636): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+640): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+644): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+648): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+652): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+656): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+660): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+664): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+668): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+672): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+676): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+680): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+684): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+688): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+692): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+696): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+700): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+704): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+708): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+712): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+716): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+720): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+724): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+728): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+732): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+736): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+740): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+744): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+748): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+752): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+756): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+760): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+764): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+768): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+772): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+776): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+780): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+784): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+788): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+792): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+796): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+800): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+804): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+808): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+812): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+816): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+820): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+824): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+828): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+832): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+836): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+840): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+844): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+848): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+852): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+856): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+860): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+864): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+868): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+872): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+876): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+880): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+884): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+888): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+892): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+896): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+900): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+904): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+908): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+912): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+916): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+920): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+924): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+928): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+932): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+936): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+940): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+944): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+948): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+952): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+956): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+960): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+964): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+968): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+972): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+976): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+980): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+984): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+988): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+992): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+996): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1000): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1004): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1008): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1012): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1016): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1020): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1024): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1028): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1032): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1036): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1040): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1044): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1048): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1052): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1056): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1060): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1064): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1068): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1072): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1076): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1080): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1084): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1088): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1092): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1096): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1100): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1104): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1108): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1112): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1116): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1120): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1124): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1128): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1132): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1136): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1140): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1144): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1148): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1152): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1156): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1160): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1164): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1168): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1172): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1176): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1180): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1184): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1188): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1192): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1196): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1200): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1204): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1208): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1212): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1216): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1220): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1224): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1228): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1232): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1236): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1240): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1244): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1248): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1252): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1256): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1260): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1264): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1268): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1272): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1276): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1280): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1284): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1288): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1292): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1296): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1300): begin 
          AHB_INTERFACE_0_hrdata<=32'h02020000; 
          end
         (32'h4000_0000+1304): begin 
          AHB_INTERFACE_0_hrdata<=32'h02020202; 
          end
         (32'h4000_0000+1308): begin 
          AHB_INTERFACE_0_hrdata<=32'h13020202; 
          end
         (32'h4000_0000+1312): begin 
          AHB_INTERFACE_0_hrdata<=32'h15151313; 
          end
         (32'h4000_0000+1316): begin 
          AHB_INTERFACE_0_hrdata<=32'h1b1b1b15; 
          end
         (32'h4000_0000+1320): begin 
          AHB_INTERFACE_0_hrdata<=32'h19040404; 
          end
         (32'h4000_0000+1324): begin 
          AHB_INTERFACE_0_hrdata<=32'h27271919; 
          end
         (32'h4000_0000+1328): begin 
          AHB_INTERFACE_0_hrdata<=32'h26262627; 
          end
         (32'h4000_0000+1332): begin 
          AHB_INTERFACE_0_hrdata<=32'h00131313; 
          end
         (32'h4000_0000+1336): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1340): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1344): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1348): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1352): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1356): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1360): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1364): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1368): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1372): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1376): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1380): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1384): begin 
          AHB_INTERFACE_0_hrdata<=32'h02020000; 
          end
         (32'h4000_0000+1388): begin 
          AHB_INTERFACE_0_hrdata<=32'h02020202; 
          end
         (32'h4000_0000+1392): begin 
          AHB_INTERFACE_0_hrdata<=32'h13020202; 
          end
         (32'h4000_0000+1396): begin 
          AHB_INTERFACE_0_hrdata<=32'h15151313; 
          end
         (32'h4000_0000+1400): begin 
          AHB_INTERFACE_0_hrdata<=32'h1b1b1b15; 
          end
         (32'h4000_0000+1404): begin 
          AHB_INTERFACE_0_hrdata<=32'h19040404; 
          end
         (32'h4000_0000+1408): begin 
          AHB_INTERFACE_0_hrdata<=32'h27271919; 
          end
         (32'h4000_0000+1412): begin 
          AHB_INTERFACE_0_hrdata<=32'h26262627; 
          end
         (32'h4000_0000+1416): begin 
          AHB_INTERFACE_0_hrdata<=32'h00131313; 
          end
         (32'h4000_0000+1420): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1424): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1428): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1432): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1436): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1440): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1444): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1448): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1452): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1456): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1460): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1464): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1468): begin 
          AHB_INTERFACE_0_hrdata<=32'h02020000; 
          end
         (32'h4000_0000+1472): begin 
          AHB_INTERFACE_0_hrdata<=32'h02020202; 
          end
         (32'h4000_0000+1476): begin 
          AHB_INTERFACE_0_hrdata<=32'h13020202; 
          end
         (32'h4000_0000+1480): begin 
          AHB_INTERFACE_0_hrdata<=32'h15151313; 
          end
         (32'h4000_0000+1484): begin 
          AHB_INTERFACE_0_hrdata<=32'h1b1b1b15; 
          end
         (32'h4000_0000+1488): begin 
          AHB_INTERFACE_0_hrdata<=32'h19040404; 
          end
         (32'h4000_0000+1492): begin 
          AHB_INTERFACE_0_hrdata<=32'h27271919; 
          end
         (32'h4000_0000+1496): begin 
          AHB_INTERFACE_0_hrdata<=32'h26262627; 
          end
         (32'h4000_0000+1500): begin 
          AHB_INTERFACE_0_hrdata<=32'h00131313; 
          end
         (32'h4000_0000+1504): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1508): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1512): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1516): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1520): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1524): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1528): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1532): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1536): begin 
          AHB_INTERFACE_0_hrdata<=32'h04000000; 
          end
         (32'h4000_0000+1540): begin 
          AHB_INTERFACE_0_hrdata<=32'h05050404; 
          end
         (32'h4000_0000+1544): begin 
          AHB_INTERFACE_0_hrdata<=32'h0e0e0e05; 
          end
         (32'h4000_0000+1548): begin 
          AHB_INTERFACE_0_hrdata<=32'h1a181818; 
          end
         (32'h4000_0000+1552): begin 
          AHB_INTERFACE_0_hrdata<=32'h27271a1a; 
          end
         (32'h4000_0000+1556): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1560): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1564): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1568): begin 
          AHB_INTERFACE_0_hrdata<=32'h23232327; 
          end
         (32'h4000_0000+1572): begin 
          AHB_INTERFACE_0_hrdata<=32'h271a1a1a; 
          end
         (32'h4000_0000+1576): begin 
          AHB_INTERFACE_0_hrdata<=32'h25252727; 
          end
         (32'h4000_0000+1580): begin 
          AHB_INTERFACE_0_hrdata<=32'h1e1e1e25; 
          end
         (32'h4000_0000+1584): begin 
          AHB_INTERFACE_0_hrdata<=32'h000a0a0a; 
          end
         (32'h4000_0000+1588): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1592): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1596): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1600): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1604): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1608): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1612): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1616): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1620): begin 
          AHB_INTERFACE_0_hrdata<=32'h04000000; 
          end
         (32'h4000_0000+1624): begin 
          AHB_INTERFACE_0_hrdata<=32'h05050404; 
          end
         (32'h4000_0000+1628): begin 
          AHB_INTERFACE_0_hrdata<=32'h0e0e0e05; 
          end
         (32'h4000_0000+1632): begin 
          AHB_INTERFACE_0_hrdata<=32'h1a181818; 
          end
         (32'h4000_0000+1636): begin 
          AHB_INTERFACE_0_hrdata<=32'h27271a1a; 
          end
         (32'h4000_0000+1640): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1644): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1648): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1652): begin 
          AHB_INTERFACE_0_hrdata<=32'h23232327; 
          end
         (32'h4000_0000+1656): begin 
          AHB_INTERFACE_0_hrdata<=32'h271a1a1a; 
          end
         (32'h4000_0000+1660): begin 
          AHB_INTERFACE_0_hrdata<=32'h25252727; 
          end
         (32'h4000_0000+1664): begin 
          AHB_INTERFACE_0_hrdata<=32'h1e1e1e25; 
          end
         (32'h4000_0000+1668): begin 
          AHB_INTERFACE_0_hrdata<=32'h000a0a0a; 
          end
         (32'h4000_0000+1672): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1676): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1680): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1684): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1688): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1692): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1696): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1700): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1704): begin 
          AHB_INTERFACE_0_hrdata<=32'h04000000; 
          end
         (32'h4000_0000+1708): begin 
          AHB_INTERFACE_0_hrdata<=32'h05050404; 
          end
         (32'h4000_0000+1712): begin 
          AHB_INTERFACE_0_hrdata<=32'h0e0e0e05; 
          end
         (32'h4000_0000+1716): begin 
          AHB_INTERFACE_0_hrdata<=32'h1a181818; 
          end
         (32'h4000_0000+1720): begin 
          AHB_INTERFACE_0_hrdata<=32'h27271a1a; 
          end
         (32'h4000_0000+1724): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1728): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1732): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1736): begin 
          AHB_INTERFACE_0_hrdata<=32'h23232327; 
          end
         (32'h4000_0000+1740): begin 
          AHB_INTERFACE_0_hrdata<=32'h271a1a1a; 
          end
         (32'h4000_0000+1744): begin 
          AHB_INTERFACE_0_hrdata<=32'h25252727; 
          end
         (32'h4000_0000+1748): begin 
          AHB_INTERFACE_0_hrdata<=32'h1e1e1e25; 
          end
         (32'h4000_0000+1752): begin 
          AHB_INTERFACE_0_hrdata<=32'h000a0a0a; 
          end
         (32'h4000_0000+1756): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1760): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1764): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1768): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1772): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1776): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1780): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1784): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1788): begin 
          AHB_INTERFACE_0_hrdata<=32'h25070707; 
          end
         (32'h4000_0000+1792): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272525; 
          end
         (32'h4000_0000+1796): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1800): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1804): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1808): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1812): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1816): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1820): begin 
          AHB_INTERFACE_0_hrdata<=32'h0e0e0e27; 
          end
         (32'h4000_0000+1824): begin 
          AHB_INTERFACE_0_hrdata<=32'h0c0c0c0c; 
          end
         (32'h4000_0000+1828): begin 
          AHB_INTERFACE_0_hrdata<=32'h08080c0c; 
          end
         (32'h4000_0000+1832): begin 
          AHB_INTERFACE_0_hrdata<=32'h05050508; 
          end
         (32'h4000_0000+1836): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1840): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1844): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1848): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1852): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1856): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1860): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1864): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1868): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1872): begin 
          AHB_INTERFACE_0_hrdata<=32'h25070707; 
          end
         (32'h4000_0000+1876): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272525; 
          end
         (32'h4000_0000+1880): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1884): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1888): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1892): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1896): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1900): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1904): begin 
          AHB_INTERFACE_0_hrdata<=32'h0e0e0e27; 
          end
         (32'h4000_0000+1908): begin 
          AHB_INTERFACE_0_hrdata<=32'h0c0c0c0c; 
          end
         (32'h4000_0000+1912): begin 
          AHB_INTERFACE_0_hrdata<=32'h08080c0c; 
          end
         (32'h4000_0000+1916): begin 
          AHB_INTERFACE_0_hrdata<=32'h05050508; 
          end
         (32'h4000_0000+1920): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1924): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1928): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1932): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1936): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1940): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1944): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1948): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1952): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+1956): begin 
          AHB_INTERFACE_0_hrdata<=32'h25070707; 
          end
         (32'h4000_0000+1960): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272525; 
          end
         (32'h4000_0000+1964): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1968): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1972): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1976): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1980): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1984): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+1988): begin 
          AHB_INTERFACE_0_hrdata<=32'h0e0e0e27; 
          end
         (32'h4000_0000+1992): begin 
          AHB_INTERFACE_0_hrdata<=32'h0c0c0c0c; 
          end
         (32'h4000_0000+1996): begin 
          AHB_INTERFACE_0_hrdata<=32'h08080c0c; 
          end
         (32'h4000_0000+2000): begin 
          AHB_INTERFACE_0_hrdata<=32'h05050508; 
          end
         (32'h4000_0000+2004): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2008): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2012): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2016): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2020): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2024): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2028): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2032): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2036): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2040): begin 
          AHB_INTERFACE_0_hrdata<=32'h22020202; 
          end
         (32'h4000_0000+2044): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272222; 
          end
         (32'h4000_0000+2048): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+2052): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+2056): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+2060): begin 
          AHB_INTERFACE_0_hrdata<=32'h1e1e1e27; 
          end
         (32'h4000_0000+2064): begin 
          AHB_INTERFACE_0_hrdata<=32'h261c1c1c; 
          end
         (32'h4000_0000+2068): begin 
          AHB_INTERFACE_0_hrdata<=32'h25252626; 
          end
         (32'h4000_0000+2072): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000025; 
          end
         (32'h4000_0000+2076): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2080): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2084): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2088): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2092): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2096): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2100): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2104): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2108): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2112): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2116): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2120): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2124): begin 
          AHB_INTERFACE_0_hrdata<=32'h22020202; 
          end
         (32'h4000_0000+2128): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272222; 
          end
         (32'h4000_0000+2132): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+2136): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+2140): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+2144): begin 
          AHB_INTERFACE_0_hrdata<=32'h1e1e1e27; 
          end
         (32'h4000_0000+2148): begin 
          AHB_INTERFACE_0_hrdata<=32'h261c1c1c; 
          end
         (32'h4000_0000+2152): begin 
          AHB_INTERFACE_0_hrdata<=32'h25252626; 
          end
         (32'h4000_0000+2156): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000025; 
          end
         (32'h4000_0000+2160): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2164): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2168): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2172): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2176): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2180): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2184): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2188): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2192): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2196): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2200): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2204): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2208): begin 
          AHB_INTERFACE_0_hrdata<=32'h22020202; 
          end
         (32'h4000_0000+2212): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272222; 
          end
         (32'h4000_0000+2216): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+2220): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+2224): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+2228): begin 
          AHB_INTERFACE_0_hrdata<=32'h1e1e1e27; 
          end
         (32'h4000_0000+2232): begin 
          AHB_INTERFACE_0_hrdata<=32'h261c1c1c; 
          end
         (32'h4000_0000+2236): begin 
          AHB_INTERFACE_0_hrdata<=32'h25252626; 
          end
         (32'h4000_0000+2240): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000025; 
          end
         (32'h4000_0000+2244): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2248): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2252): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2256): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2260): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2264): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2268): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2272): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2276): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2280): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2284): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2288): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2292): begin 
          AHB_INTERFACE_0_hrdata<=32'h0c000000; 
          end
         (32'h4000_0000+2296): begin 
          AHB_INTERFACE_0_hrdata<=32'h18180c0c; 
          end
         (32'h4000_0000+2300): begin 
          AHB_INTERFACE_0_hrdata<=32'h10101018; 
          end
         (32'h4000_0000+2304): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+2308): begin 
          AHB_INTERFACE_0_hrdata<=32'h1f1f2727; 
          end
         (32'h4000_0000+2312): begin 
          AHB_INTERFACE_0_hrdata<=32'h0101011f; 
          end
         (32'h4000_0000+2316): begin 
          AHB_INTERFACE_0_hrdata<=32'h06000000; 
          end
         (32'h4000_0000+2320): begin 
          AHB_INTERFACE_0_hrdata<=32'h18180606; 
          end
         (32'h4000_0000+2324): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000018; 
          end
         (32'h4000_0000+2328): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2332): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2336): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2340): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2344): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2348): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2352): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2356): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2360): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2364): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2368): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2372): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2376): begin 
          AHB_INTERFACE_0_hrdata<=32'h0c000000; 
          end
         (32'h4000_0000+2380): begin 
          AHB_INTERFACE_0_hrdata<=32'h18180c0c; 
          end
         (32'h4000_0000+2384): begin 
          AHB_INTERFACE_0_hrdata<=32'h10101018; 
          end
         (32'h4000_0000+2388): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+2392): begin 
          AHB_INTERFACE_0_hrdata<=32'h1f1f2727; 
          end
         (32'h4000_0000+2396): begin 
          AHB_INTERFACE_0_hrdata<=32'h0101011f; 
          end
         (32'h4000_0000+2400): begin 
          AHB_INTERFACE_0_hrdata<=32'h06000000; 
          end
         (32'h4000_0000+2404): begin 
          AHB_INTERFACE_0_hrdata<=32'h18180606; 
          end
         (32'h4000_0000+2408): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000018; 
          end
         (32'h4000_0000+2412): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2416): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2420): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2424): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2428): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2432): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2436): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2440): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2444): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2448): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2452): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2456): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2460): begin 
          AHB_INTERFACE_0_hrdata<=32'h0c000000; 
          end
         (32'h4000_0000+2464): begin 
          AHB_INTERFACE_0_hrdata<=32'h18180c0c; 
          end
         (32'h4000_0000+2468): begin 
          AHB_INTERFACE_0_hrdata<=32'h10101018; 
          end
         (32'h4000_0000+2472): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+2476): begin 
          AHB_INTERFACE_0_hrdata<=32'h1f1f2727; 
          end
         (32'h4000_0000+2480): begin 
          AHB_INTERFACE_0_hrdata<=32'h0101011f; 
          end
         (32'h4000_0000+2484): begin 
          AHB_INTERFACE_0_hrdata<=32'h06000000; 
          end
         (32'h4000_0000+2488): begin 
          AHB_INTERFACE_0_hrdata<=32'h18180606; 
          end
         (32'h4000_0000+2492): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000018; 
          end
         (32'h4000_0000+2496): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2500): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2504): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2508): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2512): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2516): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2520): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2524): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2528): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2532): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2536): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2540): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2544): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2548): begin 
          AHB_INTERFACE_0_hrdata<=32'h02020000; 
          end
         (32'h4000_0000+2552): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000002; 
          end
         (32'h4000_0000+2556): begin 
          AHB_INTERFACE_0_hrdata<=32'h27181818; 
          end
         (32'h4000_0000+2560): begin 
          AHB_INTERFACE_0_hrdata<=32'h0e0e2727; 
          end
         (32'h4000_0000+2564): begin 
          AHB_INTERFACE_0_hrdata<=32'h0000000e; 
          end
         (32'h4000_0000+2568): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2572): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2576): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2580): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2584): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2588): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2592): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2596): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2600): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2604): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2608): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2612): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2616): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2620): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2624): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2628): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2632): begin 
          AHB_INTERFACE_0_hrdata<=32'h02020000; 
          end
         (32'h4000_0000+2636): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000002; 
          end
         (32'h4000_0000+2640): begin 
          AHB_INTERFACE_0_hrdata<=32'h27181818; 
          end
         (32'h4000_0000+2644): begin 
          AHB_INTERFACE_0_hrdata<=32'h0e0e2727; 
          end
         (32'h4000_0000+2648): begin 
          AHB_INTERFACE_0_hrdata<=32'h0000000e; 
          end
         (32'h4000_0000+2652): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2656): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2660): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2664): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2668): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2672): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2676): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2680): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2684): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2688): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2692): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2696): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2700): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2704): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2708): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2712): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2716): begin 
          AHB_INTERFACE_0_hrdata<=32'h02020000; 
          end
         (32'h4000_0000+2720): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000002; 
          end
         (32'h4000_0000+2724): begin 
          AHB_INTERFACE_0_hrdata<=32'h27181818; 
          end
         (32'h4000_0000+2728): begin 
          AHB_INTERFACE_0_hrdata<=32'h0e0e2727; 
          end
         (32'h4000_0000+2732): begin 
          AHB_INTERFACE_0_hrdata<=32'h0000000e; 
          end
         (32'h4000_0000+2736): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2740): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2744): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2748): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2752): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2756): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2760): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2764): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2768): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2772): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2776): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2780): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2784): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2788): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2792): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2796): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2800): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2804): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2808): begin 
          AHB_INTERFACE_0_hrdata<=32'h27151515; 
          end
         (32'h4000_0000+2812): begin 
          AHB_INTERFACE_0_hrdata<=32'h1d1d2727; 
          end
         (32'h4000_0000+2816): begin 
          AHB_INTERFACE_0_hrdata<=32'h0000001d; 
          end
         (32'h4000_0000+2820): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2824): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2828): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2832): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2836): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2840): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2844): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2848): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2852): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2856): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2860): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2864): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2868): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2872): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2876): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2880): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2884): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2888): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2892): begin 
          AHB_INTERFACE_0_hrdata<=32'h27151515; 
          end
         (32'h4000_0000+2896): begin 
          AHB_INTERFACE_0_hrdata<=32'h1d1d2727; 
          end
         (32'h4000_0000+2900): begin 
          AHB_INTERFACE_0_hrdata<=32'h0000001d; 
          end
         (32'h4000_0000+2904): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2908): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2912): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2916): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2920): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2924): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2928): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2932): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2936): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2940): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2944): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2948): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2952): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2956): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2960): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2964): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2968): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2972): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2976): begin 
          AHB_INTERFACE_0_hrdata<=32'h27151515; 
          end
         (32'h4000_0000+2980): begin 
          AHB_INTERFACE_0_hrdata<=32'h1d1d2727; 
          end
         (32'h4000_0000+2984): begin 
          AHB_INTERFACE_0_hrdata<=32'h0000001d; 
          end
         (32'h4000_0000+2988): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2992): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+2996): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3000): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3004): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3008): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3012): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3016): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3020): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3024): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3028): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3032): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3036): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3040): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3044): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3048): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3052): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3056): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3060): begin 
          AHB_INTERFACE_0_hrdata<=32'h1d010101; 
          end
         (32'h4000_0000+3064): begin 
          AHB_INTERFACE_0_hrdata<=32'h27271d1d; 
          end
         (32'h4000_0000+3068): begin 
          AHB_INTERFACE_0_hrdata<=32'h0a0a0a27; 
          end
         (32'h4000_0000+3072): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3076): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3080): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3084): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3088): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3092): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3096): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3100): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3104): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3108): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3112): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3116): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3120): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3124): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3128): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3132): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3136): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3140): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3144): begin 
          AHB_INTERFACE_0_hrdata<=32'h1d010101; 
          end
         (32'h4000_0000+3148): begin 
          AHB_INTERFACE_0_hrdata<=32'h27271d1d; 
          end
         (32'h4000_0000+3152): begin 
          AHB_INTERFACE_0_hrdata<=32'h0a0a0a27; 
          end
         (32'h4000_0000+3156): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3160): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3164): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3168): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3172): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3176): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3180): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3184): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3188): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3192): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3196): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3200): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3204): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3208): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3212): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3216): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3220): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3224): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3228): begin 
          AHB_INTERFACE_0_hrdata<=32'h1d010101; 
          end
         (32'h4000_0000+3232): begin 
          AHB_INTERFACE_0_hrdata<=32'h27271d1d; 
          end
         (32'h4000_0000+3236): begin 
          AHB_INTERFACE_0_hrdata<=32'h0a0a0a27; 
          end
         (32'h4000_0000+3240): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3244): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3248): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3252): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3256): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3260): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3264): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3268): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3272): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3276): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3280): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3284): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3288): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3292): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3296): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3300): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3304): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3308): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3312): begin 
          AHB_INTERFACE_0_hrdata<=32'h05000000; 
          end
         (32'h4000_0000+3316): begin 
          AHB_INTERFACE_0_hrdata<=32'h25250505; 
          end
         (32'h4000_0000+3320): begin 
          AHB_INTERFACE_0_hrdata<=32'h23232325; 
          end
         (32'h4000_0000+3324): begin 
          AHB_INTERFACE_0_hrdata<=32'h10191919; 
          end
         (32'h4000_0000+3328): begin 
          AHB_INTERFACE_0_hrdata<=32'h00001010; 
          end
         (32'h4000_0000+3332): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3336): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3340): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3344): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3348): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3352): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3356): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3360): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3364): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3368): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3372): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3376): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3380): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3384): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3388): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3392): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3396): begin 
          AHB_INTERFACE_0_hrdata<=32'h05000000; 
          end
         (32'h4000_0000+3400): begin 
          AHB_INTERFACE_0_hrdata<=32'h25250505; 
          end
         (32'h4000_0000+3404): begin 
          AHB_INTERFACE_0_hrdata<=32'h23232325; 
          end
         (32'h4000_0000+3408): begin 
          AHB_INTERFACE_0_hrdata<=32'h10191919; 
          end
         (32'h4000_0000+3412): begin 
          AHB_INTERFACE_0_hrdata<=32'h00001010; 
          end
         (32'h4000_0000+3416): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3420): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3424): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3428): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3432): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3436): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3440): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3444): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3448): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3452): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3456): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3460): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3464): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3468): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3472): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3476): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3480): begin 
          AHB_INTERFACE_0_hrdata<=32'h05000000; 
          end
         (32'h4000_0000+3484): begin 
          AHB_INTERFACE_0_hrdata<=32'h25250505; 
          end
         (32'h4000_0000+3488): begin 
          AHB_INTERFACE_0_hrdata<=32'h23232325; 
          end
         (32'h4000_0000+3492): begin 
          AHB_INTERFACE_0_hrdata<=32'h10191919; 
          end
         (32'h4000_0000+3496): begin 
          AHB_INTERFACE_0_hrdata<=32'h00001010; 
          end
         (32'h4000_0000+3500): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3504): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3508): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3512): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3516): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3520): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3524): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3528): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3532): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3536): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3540): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3544): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3548): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3552): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3556): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3560): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3564): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3568): begin 
          AHB_INTERFACE_0_hrdata<=32'h0c0c0000; 
          end
         (32'h4000_0000+3572): begin 
          AHB_INTERFACE_0_hrdata<=32'h2525250c; 
          end
         (32'h4000_0000+3576): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+3580): begin 
          AHB_INTERFACE_0_hrdata<=32'h12122727; 
          end
         (32'h4000_0000+3584): begin 
          AHB_INTERFACE_0_hrdata<=32'h03030312; 
          end
         (32'h4000_0000+3588): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3592): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3596): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3600): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3604): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3608): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3612): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3616): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3620): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3624): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3628): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3632): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3636): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3640): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3644): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3648): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3652): begin 
          AHB_INTERFACE_0_hrdata<=32'h0c0c0000; 
          end
         (32'h4000_0000+3656): begin 
          AHB_INTERFACE_0_hrdata<=32'h2525250c; 
          end
         (32'h4000_0000+3660): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+3664): begin 
          AHB_INTERFACE_0_hrdata<=32'h12122727; 
          end
         (32'h4000_0000+3668): begin 
          AHB_INTERFACE_0_hrdata<=32'h03030312; 
          end
         (32'h4000_0000+3672): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3676): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3680): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3684): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3688): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3692): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3696): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3700): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3704): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3708): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3712): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3716): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3720): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3724): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3728): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3732): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3736): begin 
          AHB_INTERFACE_0_hrdata<=32'h0c0c0000; 
          end
         (32'h4000_0000+3740): begin 
          AHB_INTERFACE_0_hrdata<=32'h2525250c; 
          end
         (32'h4000_0000+3744): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+3748): begin 
          AHB_INTERFACE_0_hrdata<=32'h12122727; 
          end
         (32'h4000_0000+3752): begin 
          AHB_INTERFACE_0_hrdata<=32'h03030312; 
          end
         (32'h4000_0000+3756): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3760): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3764): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3768): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3772): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3776): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3780): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3784): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3788): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3792): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3796): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3800): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3804): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3808): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3812): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3816): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3820): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3824): begin 
          AHB_INTERFACE_0_hrdata<=32'h06060600; 
          end
         (32'h4000_0000+3828): begin 
          AHB_INTERFACE_0_hrdata<=32'h271d1d1d; 
          end
         (32'h4000_0000+3832): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+3836): begin 
          AHB_INTERFACE_0_hrdata<=32'h17171727; 
          end
         (32'h4000_0000+3840): begin 
          AHB_INTERFACE_0_hrdata<=32'h00040404; 
          end
         (32'h4000_0000+3844): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3848): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3852): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3856): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3860): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3864): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3868): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3872): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3876): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3880): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3884): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3888): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3892): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3896): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3900): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3904): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3908): begin 
          AHB_INTERFACE_0_hrdata<=32'h06060600; 
          end
         (32'h4000_0000+3912): begin 
          AHB_INTERFACE_0_hrdata<=32'h271d1d1d; 
          end
         (32'h4000_0000+3916): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+3920): begin 
          AHB_INTERFACE_0_hrdata<=32'h17171727; 
          end
         (32'h4000_0000+3924): begin 
          AHB_INTERFACE_0_hrdata<=32'h00040404; 
          end
         (32'h4000_0000+3928): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3932): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3936): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3940): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3944): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3948): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3952): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3956): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3960): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3964): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3968): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3972): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3976): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3980): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3984): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3988): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+3992): begin 
          AHB_INTERFACE_0_hrdata<=32'h06060600; 
          end
         (32'h4000_0000+3996): begin 
          AHB_INTERFACE_0_hrdata<=32'h271d1d1d; 
          end
         (32'h4000_0000+4000): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+4004): begin 
          AHB_INTERFACE_0_hrdata<=32'h17171727; 
          end
         (32'h4000_0000+4008): begin 
          AHB_INTERFACE_0_hrdata<=32'h00040404; 
          end
         (32'h4000_0000+4012): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4016): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4020): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4024): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4028): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4032): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4036): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4040): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4044): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4048): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4052): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4056): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4060): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4064): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4068): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4072): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4076): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4080): begin 
          AHB_INTERFACE_0_hrdata<=32'h0e020202; 
          end
         (32'h4000_0000+4084): begin 
          AHB_INTERFACE_0_hrdata<=32'h27270e0e; 
          end
         (32'h4000_0000+4088): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+4092): begin 
          AHB_INTERFACE_0_hrdata<=32'h001d1d1d; 
          end
         (32'h4000_0000+4096): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4100): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4104): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4108): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4112): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4116): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4120): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4124): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4128): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4132): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4136): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4140): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4144): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4148): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4152): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4156): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4160): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4164): begin 
          AHB_INTERFACE_0_hrdata<=32'h0e020202; 
          end
         (32'h4000_0000+4168): begin 
          AHB_INTERFACE_0_hrdata<=32'h27270e0e; 
          end
         (32'h4000_0000+4172): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+4176): begin 
          AHB_INTERFACE_0_hrdata<=32'h001d1d1d; 
          end
         (32'h4000_0000+4180): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4184): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4188): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4192): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4196): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4200): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4204): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4208): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4212): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4216): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4220): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4224): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4228): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4232): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4236): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4240): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4244): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4248): begin 
          AHB_INTERFACE_0_hrdata<=32'h0e020202; 
          end
         (32'h4000_0000+4252): begin 
          AHB_INTERFACE_0_hrdata<=32'h27270e0e; 
          end
         (32'h4000_0000+4256): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+4260): begin 
          AHB_INTERFACE_0_hrdata<=32'h001d1d1d; 
          end
         (32'h4000_0000+4264): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4268): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4272): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4276): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4280): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4284): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4288): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4292): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4296): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4300): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4304): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4308): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4312): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4316): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4320): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4324): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4328): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4332): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4336): begin 
          AHB_INTERFACE_0_hrdata<=32'h26260000; 
          end
         (32'h4000_0000+4340): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272726; 
          end
         (32'h4000_0000+4344): begin 
          AHB_INTERFACE_0_hrdata<=32'h0a262626; 
          end
         (32'h4000_0000+4348): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000a0a; 
          end
         (32'h4000_0000+4352): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4356): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4360): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4364): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4368): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4372): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4376): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4380): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4384): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4388): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4392): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4396): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4400): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4404): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4408): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4412): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4416): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4420): begin 
          AHB_INTERFACE_0_hrdata<=32'h26260000; 
          end
         (32'h4000_0000+4424): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272726; 
          end
         (32'h4000_0000+4428): begin 
          AHB_INTERFACE_0_hrdata<=32'h0a262626; 
          end
         (32'h4000_0000+4432): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000a0a; 
          end
         (32'h4000_0000+4436): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4440): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4444): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4448): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4452): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4456): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4460): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4464): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4468): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4472): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4476): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4480): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4484): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4488): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4492): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4496): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4500): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4504): begin 
          AHB_INTERFACE_0_hrdata<=32'h26260000; 
          end
         (32'h4000_0000+4508): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272726; 
          end
         (32'h4000_0000+4512): begin 
          AHB_INTERFACE_0_hrdata<=32'h0a262626; 
          end
         (32'h4000_0000+4516): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000a0a; 
          end
         (32'h4000_0000+4520): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4524): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4528): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4532): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4536): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4540): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4544): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4548): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4552): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4556): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4560): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4564): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4568): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4572): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4576): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4580): begin 
          AHB_INTERFACE_0_hrdata<=32'h07070700; 
          end
         (32'h4000_0000+4584): begin 
          AHB_INTERFACE_0_hrdata<=32'h1c141414; 
          end
         (32'h4000_0000+4588): begin 
          AHB_INTERFACE_0_hrdata<=32'h27271c1c; 
          end
         (32'h4000_0000+4592): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+4596): begin 
          AHB_INTERFACE_0_hrdata<=32'h00202020; 
          end
         (32'h4000_0000+4600): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4604): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4608): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4612): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4616): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4620): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4624): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4628): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4632): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4636): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4640): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4644): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4648): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4652): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4656): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4660): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4664): begin 
          AHB_INTERFACE_0_hrdata<=32'h07070700; 
          end
         (32'h4000_0000+4668): begin 
          AHB_INTERFACE_0_hrdata<=32'h1c141414; 
          end
         (32'h4000_0000+4672): begin 
          AHB_INTERFACE_0_hrdata<=32'h27271c1c; 
          end
         (32'h4000_0000+4676): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+4680): begin 
          AHB_INTERFACE_0_hrdata<=32'h00202020; 
          end
         (32'h4000_0000+4684): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4688): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4692): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4696): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4700): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4704): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4708): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4712): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4716): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4720): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4724): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4728): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4732): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4736): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4740): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4744): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4748): begin 
          AHB_INTERFACE_0_hrdata<=32'h07070700; 
          end
         (32'h4000_0000+4752): begin 
          AHB_INTERFACE_0_hrdata<=32'h1c141414; 
          end
         (32'h4000_0000+4756): begin 
          AHB_INTERFACE_0_hrdata<=32'h27271c1c; 
          end
         (32'h4000_0000+4760): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+4764): begin 
          AHB_INTERFACE_0_hrdata<=32'h00202020; 
          end
         (32'h4000_0000+4768): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4772): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4776): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4780): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4784): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4788): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4792): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4796): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4800): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4804): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4808): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4812): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4816): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4820): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4824): begin 
          AHB_INTERFACE_0_hrdata<=32'h05000000; 
          end
         (32'h4000_0000+4828): begin 
          AHB_INTERFACE_0_hrdata<=32'h17170505; 
          end
         (32'h4000_0000+4832): begin 
          AHB_INTERFACE_0_hrdata<=32'h23232317; 
          end
         (32'h4000_0000+4836): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+4840): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+4844): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+4848): begin 
          AHB_INTERFACE_0_hrdata<=32'h001c1c1c; 
          end
         (32'h4000_0000+4852): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4856): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4860): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4864): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4868): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4872): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4876): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4880): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4884): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4888): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4892): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4896): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4900): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4904): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4908): begin 
          AHB_INTERFACE_0_hrdata<=32'h05000000; 
          end
         (32'h4000_0000+4912): begin 
          AHB_INTERFACE_0_hrdata<=32'h17170505; 
          end
         (32'h4000_0000+4916): begin 
          AHB_INTERFACE_0_hrdata<=32'h23232317; 
          end
         (32'h4000_0000+4920): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+4924): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+4928): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+4932): begin 
          AHB_INTERFACE_0_hrdata<=32'h001c1c1c; 
          end
         (32'h4000_0000+4936): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4940): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4944): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4948): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4952): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4956): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4960): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4964): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4968): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4972): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4976): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4980): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4984): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4988): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+4992): begin 
          AHB_INTERFACE_0_hrdata<=32'h05000000; 
          end
         (32'h4000_0000+4996): begin 
          AHB_INTERFACE_0_hrdata<=32'h17170505; 
          end
         (32'h4000_0000+5000): begin 
          AHB_INTERFACE_0_hrdata<=32'h23232317; 
          end
         (32'h4000_0000+5004): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5008): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5012): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5016): begin 
          AHB_INTERFACE_0_hrdata<=32'h001c1c1c; 
          end
         (32'h4000_0000+5020): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5024): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5028): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5032): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5036): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5040): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5044): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5048): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5052): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5056): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5060): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5064): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5068): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5072): begin 
          AHB_INTERFACE_0_hrdata<=32'h03030300; 
          end
         (32'h4000_0000+5076): begin 
          AHB_INTERFACE_0_hrdata<=32'h22111111; 
          end
         (32'h4000_0000+5080): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272222; 
          end
         (32'h4000_0000+5084): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5088): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5092): begin 
          AHB_INTERFACE_0_hrdata<=32'h1f1f2727; 
          end
         (32'h4000_0000+5096): begin 
          AHB_INTERFACE_0_hrdata<=32'h0c0c0c1f; 
          end
         (32'h4000_0000+5100): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5104): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5108): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5112): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5116): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5120): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5124): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5128): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5132): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5136): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5140): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5144): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5148): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5152): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5156): begin 
          AHB_INTERFACE_0_hrdata<=32'h03030300; 
          end
         (32'h4000_0000+5160): begin 
          AHB_INTERFACE_0_hrdata<=32'h22111111; 
          end
         (32'h4000_0000+5164): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272222; 
          end
         (32'h4000_0000+5168): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5172): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5176): begin 
          AHB_INTERFACE_0_hrdata<=32'h1f1f2727; 
          end
         (32'h4000_0000+5180): begin 
          AHB_INTERFACE_0_hrdata<=32'h0c0c0c1f; 
          end
         (32'h4000_0000+5184): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5188): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5192): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5196): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5200): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5204): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5208): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5212): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5216): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5220): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5224): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5228): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5232): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5236): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5240): begin 
          AHB_INTERFACE_0_hrdata<=32'h03030300; 
          end
         (32'h4000_0000+5244): begin 
          AHB_INTERFACE_0_hrdata<=32'h22111111; 
          end
         (32'h4000_0000+5248): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272222; 
          end
         (32'h4000_0000+5252): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5256): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5260): begin 
          AHB_INTERFACE_0_hrdata<=32'h1f1f2727; 
          end
         (32'h4000_0000+5264): begin 
          AHB_INTERFACE_0_hrdata<=32'h0c0c0c1f; 
          end
         (32'h4000_0000+5268): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5272): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5276): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5280): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5284): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5288): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5292): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5296): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5300): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5304): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5308): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5312): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5316): begin 
          AHB_INTERFACE_0_hrdata<=32'h03000000; 
          end
         (32'h4000_0000+5320): begin 
          AHB_INTERFACE_0_hrdata<=32'h0a0a0303; 
          end
         (32'h4000_0000+5324): begin 
          AHB_INTERFACE_0_hrdata<=32'h2121210a; 
          end
         (32'h4000_0000+5328): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5332): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5336): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5340): begin 
          AHB_INTERFACE_0_hrdata<=32'h0c1e1e1e; 
          end
         (32'h4000_0000+5344): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000c0c; 
          end
         (32'h4000_0000+5348): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5352): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5356): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5360): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5364): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5368): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5372): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5376): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5380): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5384): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5388): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5392): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5396): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5400): begin 
          AHB_INTERFACE_0_hrdata<=32'h03000000; 
          end
         (32'h4000_0000+5404): begin 
          AHB_INTERFACE_0_hrdata<=32'h0a0a0303; 
          end
         (32'h4000_0000+5408): begin 
          AHB_INTERFACE_0_hrdata<=32'h2121210a; 
          end
         (32'h4000_0000+5412): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5416): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5420): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5424): begin 
          AHB_INTERFACE_0_hrdata<=32'h0c1e1e1e; 
          end
         (32'h4000_0000+5428): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000c0c; 
          end
         (32'h4000_0000+5432): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5436): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5440): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5444): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5448): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5452): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5456): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5460): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5464): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5468): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5472): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5476): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5480): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5484): begin 
          AHB_INTERFACE_0_hrdata<=32'h03000000; 
          end
         (32'h4000_0000+5488): begin 
          AHB_INTERFACE_0_hrdata<=32'h0a0a0303; 
          end
         (32'h4000_0000+5492): begin 
          AHB_INTERFACE_0_hrdata<=32'h2121210a; 
          end
         (32'h4000_0000+5496): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5500): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5504): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5508): begin 
          AHB_INTERFACE_0_hrdata<=32'h0c1e1e1e; 
          end
         (32'h4000_0000+5512): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000c0c; 
          end
         (32'h4000_0000+5516): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5520): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5524): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5528): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5532): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5536): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5540): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5544): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5548): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5552): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5556): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5560): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5564): begin 
          AHB_INTERFACE_0_hrdata<=32'h02020200; 
          end
         (32'h4000_0000+5568): begin 
          AHB_INTERFACE_0_hrdata<=32'h221a1a1a; 
          end
         (32'h4000_0000+5572): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272222; 
          end
         (32'h4000_0000+5576): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5580): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5584): begin 
          AHB_INTERFACE_0_hrdata<=32'h1e1e2727; 
          end
         (32'h4000_0000+5588): begin 
          AHB_INTERFACE_0_hrdata<=32'h0c0c0c1e; 
          end
         (32'h4000_0000+5592): begin 
          AHB_INTERFACE_0_hrdata<=32'h00010101; 
          end
         (32'h4000_0000+5596): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5600): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5604): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5608): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5612): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5616): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5620): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5624): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5628): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5632): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5636): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5640): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5644): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5648): begin 
          AHB_INTERFACE_0_hrdata<=32'h02020200; 
          end
         (32'h4000_0000+5652): begin 
          AHB_INTERFACE_0_hrdata<=32'h221a1a1a; 
          end
         (32'h4000_0000+5656): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272222; 
          end
         (32'h4000_0000+5660): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5664): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5668): begin 
          AHB_INTERFACE_0_hrdata<=32'h1e1e2727; 
          end
         (32'h4000_0000+5672): begin 
          AHB_INTERFACE_0_hrdata<=32'h0c0c0c1e; 
          end
         (32'h4000_0000+5676): begin 
          AHB_INTERFACE_0_hrdata<=32'h00010101; 
          end
         (32'h4000_0000+5680): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5684): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5688): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5692): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5696): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5700): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5704): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5708): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5712): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5716): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5720): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5724): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5728): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5732): begin 
          AHB_INTERFACE_0_hrdata<=32'h02020200; 
          end
         (32'h4000_0000+5736): begin 
          AHB_INTERFACE_0_hrdata<=32'h221a1a1a; 
          end
         (32'h4000_0000+5740): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272222; 
          end
         (32'h4000_0000+5744): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5748): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5752): begin 
          AHB_INTERFACE_0_hrdata<=32'h1e1e2727; 
          end
         (32'h4000_0000+5756): begin 
          AHB_INTERFACE_0_hrdata<=32'h0c0c0c1e; 
          end
         (32'h4000_0000+5760): begin 
          AHB_INTERFACE_0_hrdata<=32'h00010101; 
          end
         (32'h4000_0000+5764): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5768): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5772): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5776): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5780): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5784): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5788): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5792): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5796): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5800): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5804): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5808): begin 
          AHB_INTERFACE_0_hrdata<=32'h08000000; 
          end
         (32'h4000_0000+5812): begin 
          AHB_INTERFACE_0_hrdata<=32'h1a1a0808; 
          end
         (32'h4000_0000+5816): begin 
          AHB_INTERFACE_0_hrdata<=32'h2323231a; 
          end
         (32'h4000_0000+5820): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5824): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5828): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5832): begin 
          AHB_INTERFACE_0_hrdata<=32'h14262626; 
          end
         (32'h4000_0000+5836): begin 
          AHB_INTERFACE_0_hrdata<=32'h01011414; 
          end
         (32'h4000_0000+5840): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000001; 
          end
         (32'h4000_0000+5844): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5848): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5852): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5856): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5860): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5864): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5868): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5872): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5876): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5880): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5884): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5888): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5892): begin 
          AHB_INTERFACE_0_hrdata<=32'h08000000; 
          end
         (32'h4000_0000+5896): begin 
          AHB_INTERFACE_0_hrdata<=32'h1a1a0808; 
          end
         (32'h4000_0000+5900): begin 
          AHB_INTERFACE_0_hrdata<=32'h2323231a; 
          end
         (32'h4000_0000+5904): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5908): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5912): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5916): begin 
          AHB_INTERFACE_0_hrdata<=32'h14262626; 
          end
         (32'h4000_0000+5920): begin 
          AHB_INTERFACE_0_hrdata<=32'h01011414; 
          end
         (32'h4000_0000+5924): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000001; 
          end
         (32'h4000_0000+5928): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5932): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5936): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5940): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5944): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5948): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5952): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5956): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5960): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5964): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5968): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5972): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+5976): begin 
          AHB_INTERFACE_0_hrdata<=32'h08000000; 
          end
         (32'h4000_0000+5980): begin 
          AHB_INTERFACE_0_hrdata<=32'h1a1a0808; 
          end
         (32'h4000_0000+5984): begin 
          AHB_INTERFACE_0_hrdata<=32'h2323231a; 
          end
         (32'h4000_0000+5988): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5992): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+5996): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+6000): begin 
          AHB_INTERFACE_0_hrdata<=32'h14262626; 
          end
         (32'h4000_0000+6004): begin 
          AHB_INTERFACE_0_hrdata<=32'h01011414; 
          end
         (32'h4000_0000+6008): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000001; 
          end
         (32'h4000_0000+6012): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6016): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6020): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6024): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6028): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6032): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6036): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6040): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6044): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6048): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6052): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6056): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6060): begin 
          AHB_INTERFACE_0_hrdata<=32'h15000000; 
          end
         (32'h4000_0000+6064): begin 
          AHB_INTERFACE_0_hrdata<=32'h27271515; 
          end
         (32'h4000_0000+6068): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+6072): begin 
          AHB_INTERFACE_0_hrdata<=32'h21272727; 
          end
         (32'h4000_0000+6076): begin 
          AHB_INTERFACE_0_hrdata<=32'h14142121; 
          end
         (32'h4000_0000+6080): begin 
          AHB_INTERFACE_0_hrdata<=32'h14141414; 
          end
         (32'h4000_0000+6084): begin 
          AHB_INTERFACE_0_hrdata<=32'h00020202; 
          end
         (32'h4000_0000+6088): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6092): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6096): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6100): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6104): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6108): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6112): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6116): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6120): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6124): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6128): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6132): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6136): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6140): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6144): begin 
          AHB_INTERFACE_0_hrdata<=32'h15000000; 
          end
         (32'h4000_0000+6148): begin 
          AHB_INTERFACE_0_hrdata<=32'h27271515; 
          end
         (32'h4000_0000+6152): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+6156): begin 
          AHB_INTERFACE_0_hrdata<=32'h21272727; 
          end
         (32'h4000_0000+6160): begin 
          AHB_INTERFACE_0_hrdata<=32'h14142121; 
          end
         (32'h4000_0000+6164): begin 
          AHB_INTERFACE_0_hrdata<=32'h14141414; 
          end
         (32'h4000_0000+6168): begin 
          AHB_INTERFACE_0_hrdata<=32'h00020202; 
          end
         (32'h4000_0000+6172): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6176): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6180): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6184): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6188): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6192): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6196): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6200): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6204): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6208): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6212): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6216): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6220): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6224): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6228): begin 
          AHB_INTERFACE_0_hrdata<=32'h15000000; 
          end
         (32'h4000_0000+6232): begin 
          AHB_INTERFACE_0_hrdata<=32'h27271515; 
          end
         (32'h4000_0000+6236): begin 
          AHB_INTERFACE_0_hrdata<=32'h27272727; 
          end
         (32'h4000_0000+6240): begin 
          AHB_INTERFACE_0_hrdata<=32'h21272727; 
          end
         (32'h4000_0000+6244): begin 
          AHB_INTERFACE_0_hrdata<=32'h14142121; 
          end
         (32'h4000_0000+6248): begin 
          AHB_INTERFACE_0_hrdata<=32'h14141414; 
          end
         (32'h4000_0000+6252): begin 
          AHB_INTERFACE_0_hrdata<=32'h00020202; 
          end
         (32'h4000_0000+6256): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6260): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6264): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6268): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6272): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6276): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6280): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6284): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6288): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6292): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6296): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6300): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6304): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6308): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6312): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6316): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6320): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6324): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6328): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6332): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6336): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6340): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6344): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6348): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6352): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6356): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6360): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6364): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6368): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6372): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6376): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6380): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6384): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6388): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6392): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6396): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6400): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6404): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6408): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6412): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6416): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6420): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6424): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6428): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6432): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6436): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6440): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6444): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6448): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6452): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6456): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6460): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6464): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6468): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6472): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6476): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6480): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6484): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6488): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6492): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6496): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6500): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6504): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6508): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6512): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6516): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6520): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6524): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6528): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6532): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6536): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6540): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6544): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6548): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6552): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6556): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6560): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6564): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6568): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6572): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6576): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6580): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6584): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6588): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6592): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6596): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6600): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6604): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6608): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6612): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6616): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6620): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6624): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6628): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6632): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6636): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6640): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6644): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6648): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6652): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6656): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6660): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6664): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6668): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6672): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6676): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6680): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6684): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6688): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6692): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6696): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6700): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6704): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6708): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6712): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6716): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6720): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6724): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6728): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6732): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6736): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6740): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6744): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6748): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6752): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6756): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6760): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6764): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6768): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6772): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6776): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6780): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6784): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6788): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6792): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end
         (32'h4000_0000+6796): begin 
          AHB_INTERFACE_0_hrdata<=32'h00000000; 
          end

         endcase
      end
endmodule
 
